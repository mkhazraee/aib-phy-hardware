// SPDX-License-Identifier: Apache-2.0
// Copyright (C) 2019 Intel Corporation. 
//------------------------------------------------------------------------
// Copyright (c) 2012 Altera Corporation. .
// Library - aibndaux_lib, Cell - aibndaux_pasred, View - schematic
// LAST TIME SAVED: Jul  8 18:04:04 2015
// NETLIST TIME: Jul  9 10:28:17 2015
// `timescale 1ps/1ps

module aibndaux_pasred ( crete_detect, jtr_tck, jtr_tdo, jtr_tms, iopad_crdet,
     iopad_dn_por, iopad_dn_rst_n, iopad_jt_tck, iopad_jt_tdi,
     iopad_jt_tms, iopad_jtr_tck, iopad_jtr_tdo, iopad_jtr_tms,
     anlg_rstb, csr_iocsr_sel, csr_pred_dataselb, csr_pred_ndrv,
     csr_pred_pdrv, csr_pred_rxen, csr_pred_txen, dig_rstb, dn_por,
     dn_rst_n, jt_tck, jt_tdi, jt_tms, vccl_aibndaux, vssl_aibndaux );

output  crete_detect, jtr_tck, jtr_tdo, jtr_tms;

inout  iopad_crdet, iopad_dn_por, iopad_dn_rst_n, iopad_jt_tck,
     iopad_jt_tdi, iopad_jt_tms, iopad_jtr_tck, iopad_jtr_tdo,
     iopad_jtr_tms;

input  anlg_rstb, csr_iocsr_sel, csr_pred_dataselb, csr_pred_txen,
     dig_rstb, dn_por, dn_rst_n, jt_tck, jt_tdi, jt_tms, vccl_aibndaux,
     vssl_aibndaux;

input [1:0]  csr_pred_ndrv;
input [1:0]  csr_pred_pdrv;
input [2:0]  csr_pred_rxen;

wire jtr_tck, crete_detect, jtr_tck_int, jt_tck, jtr_tms, jtr_tms_int, jt_tms, jtr_tdo, jtr_tdo_int, jt_tdi, csr_iocsr_sel, vssl_aibndaux, csr_pred_txen_int, csr_pred_txen, vccl_aibndaux; // Conversion Sript Generated

// Buses in the design

wire  [2:0]  csr_pred_rxen_int;

wire  [1:0]  csr_pred_ndrv_int;

wire  [1:0]  csr_pred_pdrv_int;


// specify 
//     specparam CDS_LIBNAME  = "aibndaux_lib";
//     specparam CDS_CELLNAME = "aibndaux_pasred";
//     specparam CDS_VIEWNAME = "schematic";
// endspecify

aibnd_buffx1_top  xcrdet ( .idata1_in1_jtag_out(net0282),
     .async_dat_in1_jtag_out(net0266), .idata0_in1_jtag_out(net0310),
     .prev_io_shift_en(vssl_aibndaux), .jtag_clkdr_outn(net0203),
     .anlg_rstb(vccl_aibndaux), .pd_data_aib(net087),
     .oclk_out(net075), .oclkb_out(net076), .odat0_out(net077),
     .odat1_out(net078), .odat_async_out(crete_detect),
     .pd_data_out(net080), .async_dat_in0(vssl_aibndaux),
     .async_dat_in1(vssl_aibndaux), .iclkin_dist_in0(vssl_aibndaux),
     .iclkin_dist_in1(vssl_aibndaux), .idata0_in0(vssl_aibndaux),
     .idata0_in1(vssl_aibndaux), .idata1_in0(vssl_aibndaux),
     .idata1_in1(vssl_aibndaux), .idataselb_in0(vssl_aibndaux),
     .idataselb_in1(vssl_aibndaux), .iddren_in0(vssl_aibndaux),
     .iddren_in1(vssl_aibndaux), .ilaunch_clk_in0(vssl_aibndaux),
     .ilaunch_clk_in1(vssl_aibndaux), .ilpbk_dat_in0(vssl_aibndaux),
     .ilpbk_dat_in1(vssl_aibndaux), .ilpbk_en_in0(vssl_aibndaux),
     .ilpbk_en_in1(vssl_aibndaux), .indrv_in0({vssl_aibndaux,
     vssl_aibndaux}), .indrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .irxen_in0({vssl_aibndaux,vssl_aibndaux,vssl_aibndaux}),
     .irxen_in1({vssl_aibndaux,vssl_aibndaux,vssl_aibndaux}), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(vssl_aibndaux),
     .itxen_in1(vssl_aibndaux), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(net086), .oclkb_in1(vssl_aibndaux),
     .jtag_clksel(vssl_aibndaux), .odat0_in1(vssl_aibndaux),
     .vssl_aibnd(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(vssl_aibndaux), .shift_en(vssl_aibndaux),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net040), .jtag_intest(vssl_aibndaux),
     .odat1_aib(net085), .jtag_rx_scan_out(net041), .odat0_aib(net084),
     .oclk_aib(net082), .last_bs_out(net042),
     .vccl_aibnd(vccl_aibndaux), .oclkb_aib(net083),
     .jtag_clkdr_in(vssl_aibndaux), .jtag_rstb_en(vssl_aibndaux),
     .jtag_mode_in(vssl_aibndaux), .jtag_rstb(vssl_aibndaux),
     .jtag_tx_scan_in(vssl_aibndaux),
     .jtag_tx_scanen_in(vssl_aibndaux), .last_bs_in(vssl_aibndaux),
     .iopad(iopad_crdet), .oclkn(net081), .iclkn(vssl_aibndaux),
     .test_weakpu(vssl_aibndaux), .test_weakpd(vccl_aibndaux));
aibnd_buffx1_top  xtstmx2 ( .idata1_in1_jtag_out(net0285),
     .async_dat_in1_jtag_out(net0102), .idata0_in1_jtag_out(net0312),
     .prev_io_shift_en(vssl_aibndaux), .jtag_clkdr_outn(net0271),
     .jtag_clksel(vssl_aibndaux), .vssl_aibnd(vssl_aibndaux),
     .jtag_intest(vssl_aibndaux), .vccl_aibnd(vccl_aibndaux),
     .jtag_rstb_en(vssl_aibndaux), .anlg_rstb(anlg_rstb),
     .pd_data_aib(net0255), .oclk_out(net0206), .oclkb_out(net0210),
     .odat0_out(net0214), .odat1_out(net0218),
     .odat_async_out(jtr_tms_int), .pd_data_out(net0222),
     .async_dat_in0(vssl_aibndaux), .async_dat_in1(vssl_aibndaux),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(vssl_aibndaux), .idataselb_in1(vssl_aibndaux),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .indrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .irxen_in0(csr_pred_rxen_int[2:0]),
     .irxen_in1(csr_pred_rxen_int[2:0]), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(vssl_aibndaux),
     .itxen_in1(vssl_aibndaux), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(net0251), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(vssl_aibndaux), .shift_en(vssl_aibndaux),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net043), .odat1_aib(net0247),
     .jtag_rx_scan_out(net044), .odat0_aib(net0243),
     .oclk_aib(net0235), .last_bs_out(net045), .oclkb_aib(net0239),
     .jtag_clkdr_in(vssl_aibndaux), .jtag_mode_in(vssl_aibndaux),
     .jtag_rstb(vssl_aibndaux), .jtag_tx_scan_in(vssl_aibndaux),
     .jtag_tx_scanen_in(vssl_aibndaux), .last_bs_in(vssl_aibndaux),
     .iopad(iopad_jtr_tms), .oclkn(net0231), .iclkn(vssl_aibndaux),
     .test_weakpu(vssl_aibndaux), .test_weakpd(vssl_aibndaux));
aibnd_buffx1_top  xjt_tms ( .idata1_in1_jtag_out(net0324),
     .async_dat_in1_jtag_out(net0321), .idata0_in1_jtag_out(net094),
     .prev_io_shift_en(vssl_aibndaux), .jtag_clkdr_outn(net0284),
     .jtag_clksel(vssl_aibndaux), .vssl_aibnd(vssl_aibndaux),
     .jtag_intest(vssl_aibndaux), .vccl_aibnd(vccl_aibndaux),
     .jtag_rstb_en(vssl_aibndaux), .anlg_rstb(anlg_rstb),
     .pd_data_aib(net0253), .oclk_out(net0204), .oclkb_out(net0208),
     .odat0_out(net0212), .odat1_out(net0216),
     .odat_async_out(net0199), .pd_data_out(net0220),
     .async_dat_in0(jt_tms), .async_dat_in1(vssl_aibndaux),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(csr_pred_dataselb), .idataselb_in1(vssl_aibndaux),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0(csr_pred_ndrv_int[1:0]),
     .indrv_in1(csr_pred_ndrv_int[1:0]),
     .ipdrv_in0(csr_pred_pdrv_int[1:0]),
     .ipdrv_in1(csr_pred_pdrv_int[1:0]), .irxen_in0({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .irxen_in1({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(csr_pred_txen_int),
     .itxen_in1(csr_pred_txen_int), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(net0249), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(vssl_aibndaux), .shift_en(vssl_aibndaux),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net052), .odat1_aib(net0245),
     .jtag_rx_scan_out(net053), .odat0_aib(net0241),
     .oclk_aib(net0233), .last_bs_out(net054), .oclkb_aib(net0237),
     .jtag_clkdr_in(vssl_aibndaux), .jtag_mode_in(vssl_aibndaux),
     .jtag_rstb(vssl_aibndaux), .jtag_tx_scan_in(vssl_aibndaux),
     .jtag_tx_scanen_in(vssl_aibndaux), .last_bs_in(vssl_aibndaux),
     .iopad(iopad_jt_tms), .oclkn(net0229), .iclkn(vssl_aibndaux),
     .test_weakpu(vssl_aibndaux), .test_weakpd(vssl_aibndaux));
aibnd_buffx1_top  xjt_tdi ( .idata1_in1_jtag_out(net0275),
     .async_dat_in1_jtag_out(net0311), .idata0_in1_jtag_out(net0268),
     .prev_io_shift_en(vssl_aibndaux), .jtag_clkdr_outn(net0277),
     .jtag_clksel(vssl_aibndaux), .vssl_aibnd(vssl_aibndaux),
     .jtag_intest(vssl_aibndaux), .vccl_aibnd(vccl_aibndaux),
     .jtag_rstb_en(vssl_aibndaux), .anlg_rstb(anlg_rstb),
     .pd_data_aib(net0101), .oclk_out(net088), .oclkb_out(net089),
     .odat0_out(net090), .odat1_out(net091), .odat_async_out(net092),
     .pd_data_out(net093), .async_dat_in0(jt_tdi),
     .async_dat_in1(vssl_aibndaux), .iclkin_dist_in0(vssl_aibndaux),
     .iclkin_dist_in1(vssl_aibndaux), .idata0_in0(vssl_aibndaux),
     .idata0_in1(vssl_aibndaux), .idata1_in0(vssl_aibndaux),
     .idata1_in1(vssl_aibndaux), .idataselb_in0(csr_pred_dataselb),
     .idataselb_in1(vssl_aibndaux), .iddren_in0(vssl_aibndaux),
     .iddren_in1(vssl_aibndaux), .ilaunch_clk_in0(vssl_aibndaux),
     .ilaunch_clk_in1(vssl_aibndaux), .ilpbk_dat_in0(vssl_aibndaux),
     .ilpbk_dat_in1(vssl_aibndaux), .ilpbk_en_in0(vssl_aibndaux),
     .ilpbk_en_in1(vssl_aibndaux), .indrv_in0(csr_pred_ndrv_int[1:0]),
     .indrv_in1(csr_pred_ndrv_int[1:0]),
     .ipdrv_in0(csr_pred_pdrv_int[1:0]),
     .ipdrv_in1(csr_pred_pdrv_int[1:0]), .irxen_in0({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .irxen_in1({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(csr_pred_txen_int),
     .itxen_in1(csr_pred_txen_int), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(net0100), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(vssl_aibndaux), .shift_en(vssl_aibndaux),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net059), .odat1_aib(net099),
     .jtag_rx_scan_out(net058), .odat0_aib(net098), .oclk_aib(net096),
     .last_bs_out(net060), .oclkb_aib(net097),
     .jtag_clkdr_in(vssl_aibndaux), .jtag_mode_in(vssl_aibndaux),
     .jtag_rstb(vssl_aibndaux), .jtag_tx_scan_in(vssl_aibndaux),
     .jtag_tx_scanen_in(vssl_aibndaux), .last_bs_in(vssl_aibndaux),
     .iopad(iopad_jt_tdi), .oclkn(net095), .iclkn(vssl_aibndaux),
     .test_weakpu(vssl_aibndaux), .test_weakpd(vssl_aibndaux));
aibnd_buffx1_top  xjt_tck ( .idata1_in1_jtag_out(net0317),
     .async_dat_in1_jtag_out(net0320), .idata0_in1_jtag_out(net0287),
     .prev_io_shift_en(vssl_aibndaux), .jtag_clkdr_outn(net0274),
     .jtag_clksel(vssl_aibndaux), .vssl_aibnd(vssl_aibndaux),
     .jtag_intest(vssl_aibndaux), .vccl_aibnd(vccl_aibndaux),
     .jtag_rstb_en(vssl_aibndaux), .anlg_rstb(anlg_rstb),
     .pd_data_aib(net0263), .oclk_out(net0224), .oclkb_out(net0225),
     .odat0_out(net0226), .odat1_out(net0227),
     .odat_async_out(net0267), .pd_data_out(net0228),
     .async_dat_in0(jt_tck), .async_dat_in1(vssl_aibndaux),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(csr_pred_dataselb), .idataselb_in1(vssl_aibndaux),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0(csr_pred_ndrv_int[1:0]),
     .indrv_in1(csr_pred_ndrv_int[1:0]),
     .ipdrv_in0(csr_pred_pdrv_int[1:0]),
     .ipdrv_in1(csr_pred_pdrv_int[1:0]), .irxen_in0({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .irxen_in1({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(csr_pred_txen_int),
     .itxen_in1(csr_pred_txen_int), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(net0262), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(vssl_aibndaux), .shift_en(vssl_aibndaux),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net056), .odat1_aib(net0261),
     .jtag_rx_scan_out(net057), .odat0_aib(net0260),
     .oclk_aib(net0258), .last_bs_out(net055), .oclkb_aib(net0259),
     .jtag_clkdr_in(vssl_aibndaux), .jtag_mode_in(vssl_aibndaux),
     .jtag_rstb(vssl_aibndaux), .jtag_tx_scan_in(vssl_aibndaux),
     .jtag_tx_scanen_in(vssl_aibndaux), .last_bs_in(vssl_aibndaux),
     .iopad(iopad_jt_tck), .oclkn(net0257), .iclkn(vssl_aibndaux),
     .test_weakpu(vssl_aibndaux), .test_weakpd(vssl_aibndaux));
aibnd_buffx1_top  xdn_por ( .idata1_in1_jtag_out(net0309),
     .async_dat_in1_jtag_out(net0283), .idata0_in1_jtag_out(net0313),
     .prev_io_shift_en(vssl_aibndaux), .jtag_clkdr_outn(net0264),
     .jtag_clksel(vssl_aibndaux), .vssl_aibnd(vssl_aibndaux),
     .jtag_intest(vssl_aibndaux), .vccl_aibnd(vccl_aibndaux),
     .jtag_rstb_en(vssl_aibndaux), .anlg_rstb(vccl_aibndaux),
     .pd_data_aib(net0115), .oclk_out(net0103), .oclkb_out(net0104),
     .odat0_out(net0105), .odat1_out(net0106),
     .odat_async_out(net0107), .pd_data_out(net0108),
     .async_dat_in0(dn_por), .async_dat_in1(vssl_aibndaux),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(vssl_aibndaux), .idataselb_in1(vssl_aibndaux),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0({vccl_aibndaux, vssl_aibndaux}),
     .indrv_in1({vccl_aibndaux, vssl_aibndaux}),
     .ipdrv_in0({vccl_aibndaux, vssl_aibndaux}),
     .ipdrv_in1({vccl_aibndaux, vssl_aibndaux}), .irxen_in0({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .irxen_in1({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(csr_pred_txen_int),
     .itxen_in1(csr_pred_txen_int), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(net0114), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(vssl_aibndaux), .shift_en(vssl_aibndaux),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net061), .odat1_aib(net0113),
     .jtag_rx_scan_out(net062), .odat0_aib(net0112),
     .oclk_aib(net0110), .last_bs_out(net063), .oclkb_aib(net0111),
     .jtag_clkdr_in(vssl_aibndaux), .jtag_mode_in(vssl_aibndaux),
     .jtag_rstb(vssl_aibndaux), .jtag_tx_scan_in(vssl_aibndaux),
     .jtag_tx_scanen_in(vssl_aibndaux), .last_bs_in(vssl_aibndaux),
     .iopad(iopad_dn_por), .oclkn(net0109), .iclkn(vssl_aibndaux),
     .test_weakpu(vssl_aibndaux), .test_weakpd(vssl_aibndaux));
aibnd_buffx1_top  xdn_rst_n ( .idata1_in1_jtag_out(net0290),
     .async_dat_in1_jtag_out(net0280), .idata0_in1_jtag_out(net0307),
     .prev_io_shift_en(vssl_aibndaux), .jtag_clkdr_outn(net0278),
     .jtag_clksel(vssl_aibndaux), .vssl_aibnd(vssl_aibndaux),
     .jtag_intest(vssl_aibndaux), .vccl_aibnd(vccl_aibndaux),
     .jtag_rstb_en(vssl_aibndaux), .anlg_rstb(anlg_rstb),
     .pd_data_aib(net0130), .oclk_out(net0442), .oclkb_out(net0416),
     .odat0_out(net028), .odat1_out(net029), .odat_async_out(net0385),
     .pd_data_out(net0402), .async_dat_in0(dn_rst_n),
     .async_dat_in1(vssl_aibndaux), .iclkin_dist_in0(vssl_aibndaux),
     .iclkin_dist_in1(vssl_aibndaux), .idata0_in0(vssl_aibndaux),
     .idata0_in1(vssl_aibndaux), .idata1_in0(vssl_aibndaux),
     .idata1_in1(vssl_aibndaux), .idataselb_in0(csr_pred_dataselb),
     .idataselb_in1(vssl_aibndaux), .iddren_in0(vssl_aibndaux),
     .iddren_in1(vssl_aibndaux), .ilaunch_clk_in0(vssl_aibndaux),
     .ilaunch_clk_in1(vssl_aibndaux), .ilpbk_dat_in0(vssl_aibndaux),
     .ilpbk_dat_in1(vssl_aibndaux), .ilpbk_en_in0(vssl_aibndaux),
     .ilpbk_en_in1(vssl_aibndaux), .indrv_in0(csr_pred_ndrv_int[1:0]),
     .indrv_in1(csr_pred_ndrv_int[1:0]),
     .ipdrv_in0(csr_pred_pdrv_int[1:0]),
     .ipdrv_in1(csr_pred_pdrv_int[1:0]), .irxen_in0({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .irxen_in1({vssl_aibndaux,
     vccl_aibndaux, vssl_aibndaux}), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(csr_pred_txen_int),
     .itxen_in1(csr_pred_txen_int), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(net0129), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(vssl_aibndaux), .shift_en(vssl_aibndaux),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net066), .odat1_aib(net0128),
     .jtag_rx_scan_out(net065), .odat0_aib(net0127),
     .oclk_aib(net0125), .last_bs_out(net064), .oclkb_aib(net0126),
     .jtag_clkdr_in(vssl_aibndaux), .jtag_mode_in(vssl_aibndaux),
     .jtag_rstb(vssl_aibndaux), .jtag_tx_scan_in(vssl_aibndaux),
     .jtag_tx_scanen_in(vssl_aibndaux), .last_bs_in(vssl_aibndaux),
     .iopad(iopad_dn_rst_n), .oclkn(net0124), .iclkn(vssl_aibndaux),
     .test_weakpu(vssl_aibndaux), .test_weakpd(vssl_aibndaux));
aibnd_buffx1_top  xtstmx0 ( .idata1_in1_jtag_out(net0304),
     .async_dat_in1_jtag_out(net0323), .idata0_in1_jtag_out(net0322),
     .prev_io_shift_en(vssl_aibndaux), .jtag_clkdr_outn(net0276),
     .jtag_clksel(vssl_aibndaux), .vssl_aibnd(vssl_aibndaux),
     .jtag_intest(vssl_aibndaux), .vccl_aibnd(vccl_aibndaux),
     .jtag_rstb_en(vssl_aibndaux), .anlg_rstb(anlg_rstb),
     .pd_data_aib(net0254), .oclk_out(net0205), .oclkb_out(net0209),
     .odat0_out(net0213), .odat1_out(net0217),
     .odat_async_out(jtr_tdo_int), .pd_data_out(net0221),
     .async_dat_in0(vssl_aibndaux), .async_dat_in1(vssl_aibndaux),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(vssl_aibndaux), .idataselb_in1(vssl_aibndaux),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .indrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .irxen_in0(csr_pred_rxen_int[2:0]),
     .irxen_in1(csr_pred_rxen_int[2:0]), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(vssl_aibndaux),
     .itxen_in1(vssl_aibndaux), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(net0250), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(vssl_aibndaux), .shift_en(vssl_aibndaux),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net046), .odat1_aib(net0246),
     .jtag_rx_scan_out(net047), .odat0_aib(net0242),
     .oclk_aib(net0234), .last_bs_out(net048), .oclkb_aib(net0238),
     .jtag_clkdr_in(vssl_aibndaux), .jtag_mode_in(vssl_aibndaux),
     .jtag_rstb(vssl_aibndaux), .jtag_tx_scan_in(vssl_aibndaux),
     .jtag_tx_scanen_in(vssl_aibndaux), .last_bs_in(vssl_aibndaux),
     .iopad(iopad_jtr_tdo), .oclkn(net0230), .iclkn(vssl_aibndaux),
     .test_weakpu(vssl_aibndaux), .test_weakpd(vssl_aibndaux));
aibnd_buffx1_top  xio_oe0 ( .idata1_in1_jtag_out(net0305),
     .async_dat_in1_jtag_out(net0292), .idata0_in1_jtag_out(net0318),
     .prev_io_shift_en(vssl_aibndaux), .jtag_clkdr_outn(net0281),
     .jtag_clksel(vssl_aibndaux), .vssl_aibnd(vssl_aibndaux),
     .jtag_intest(vssl_aibndaux), .vccl_aibnd(vccl_aibndaux),
     .jtag_rstb_en(vssl_aibndaux), .anlg_rstb(anlg_rstb),
     .pd_data_aib(net0256), .oclk_out(net0207), .oclkb_out(net0211),
     .odat0_out(net0215), .odat1_out(net0219),
     .odat_async_out(jtr_tck_int), .pd_data_out(net0223),
     .async_dat_in0(vssl_aibndaux), .async_dat_in1(vssl_aibndaux),
     .iclkin_dist_in0(vssl_aibndaux), .iclkin_dist_in1(vssl_aibndaux),
     .idata0_in0(vssl_aibndaux), .idata0_in1(vssl_aibndaux),
     .idata1_in0(vssl_aibndaux), .idata1_in1(vssl_aibndaux),
     .idataselb_in0(vssl_aibndaux), .idataselb_in1(vssl_aibndaux),
     .iddren_in0(vssl_aibndaux), .iddren_in1(vssl_aibndaux),
     .ilaunch_clk_in0(vssl_aibndaux), .ilaunch_clk_in1(vssl_aibndaux),
     .ilpbk_dat_in0(vssl_aibndaux), .ilpbk_dat_in1(vssl_aibndaux),
     .ilpbk_en_in0(vssl_aibndaux), .ilpbk_en_in1(vssl_aibndaux),
     .indrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .indrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in0({vssl_aibndaux, vssl_aibndaux}),
     .ipdrv_in1({vssl_aibndaux, vssl_aibndaux}),
     .irxen_in0(csr_pred_rxen_int[2:0]),
     .irxen_in1(csr_pred_rxen_int[2:0]), .istrbclk_in0(vssl_aibndaux),
     .istrbclk_in1(vssl_aibndaux), .itxen_in0(vssl_aibndaux),
     .itxen_in1(vssl_aibndaux), .oclk_in1(vssl_aibndaux),
     .odat_async_aib(net0252), .oclkb_in1(vssl_aibndaux),
     .odat0_in1(vssl_aibndaux), .odat1_in1(vssl_aibndaux),
     .odat_async_in1(vssl_aibndaux), .shift_en(vssl_aibndaux),
     .pd_data_in1(vssl_aibndaux), .dig_rstb(dig_rstb),
     .jtag_clkdr_out(net051), .odat1_aib(net0248),
     .jtag_rx_scan_out(net050), .odat0_aib(net0244),
     .oclk_aib(net0236), .last_bs_out(net049), .oclkb_aib(net0240),
     .jtag_clkdr_in(vssl_aibndaux), .jtag_mode_in(vssl_aibndaux),
     .jtag_rstb(vssl_aibndaux), .jtag_tx_scan_in(vssl_aibndaux),
     .jtag_tx_scanen_in(vssl_aibndaux), .last_bs_in(vssl_aibndaux),
     .iopad(iopad_jtr_tck), .oclkn(net0232), .iclkn(vssl_aibndaux),
     .test_weakpu(vssl_aibndaux), .test_weakpd(vssl_aibndaux));

assign jtr_tck = crete_detect ? jtr_tck_int : jt_tck;
assign jtr_tms = crete_detect ? jtr_tms_int : jt_tms;
assign jtr_tdo = crete_detect ? jtr_tdo_int : jt_tdi;
assign csr_pred_ndrv_int[1:0] = csr_iocsr_sel ? csr_pred_ndrv[1:0] : {vccl_aibndaux, vssl_aibndaux};
assign csr_pred_pdrv_int[1:0] = csr_iocsr_sel ? csr_pred_pdrv[1:0] : {vccl_aibndaux, vssl_aibndaux};
assign csr_pred_rxen_int[2:0] = csr_iocsr_sel ? csr_pred_rxen[2:0] : vssl_aibndaux;
assign csr_pred_txen_int = csr_iocsr_sel ? csr_pred_txen : crete_detect;


endmodule

