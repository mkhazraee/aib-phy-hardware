// SPDX-License-Identifier: Apache-2.0
// Copyright (C) 2019 Intel Corporation. 
// Library - aibnd_lib, Cell - aibnd_avmm1, View - schematic
// LAST TIME SAVED: Jul  6 22:41:38 2015
// NETLIST TIME: Jul  8 13:09:51 2015
// `timescale 1ps/1ps

module aibnd_avmm1 ( avmm1_odat0, avmm1_odat1, avmm2_rx_distclk,
     avmm2_rx_strbclk, avmm2_tx_launch_clk_l0, avmm2_tx_launch_clk_l1,
     iclkin_dist_vinp0, iclkin_dist_vinp1, idat0_voutp00,
     idat0_voutp01, idat1_voutp00, idat1_voutp01, idata0_ssrdout,
     idata0_ssrldout, idata1_ssrdout, idata1_ssrldout,
     idataselb_ssrdout, idataselb_ssrldout, idataselb_voutp00,
     idataselb_voutp01, ilaunch_clk_ssrdout, ilaunch_clk_ssrldout,
     ilaunch_clk_voutp00, ilaunch_clk_voutp01, irxen_vinp0,
     istrbclk_vinp0, istrbclk_vinp1, itxen_ssrdout, itxen_ssrldout,
     itxen_voutp00, itxen_voutp01, jtag_clkdr_in_srcclkinn,
     jtag_clkdr_in_ssrdout, jtag_clkdr_in_ssrldout, jtag_clkdr_vinp0,
     jtag_clkdr_voutp00, jtag_clkdr_voutp01, jtag_rx_scan_in_srcclkinn,
     jtag_rx_scan_in_ssrdout, jtag_rx_scan_in_ssrldout,
     jtag_rx_scan_vinp0, jtag_rx_scan_voutp00, jtag_rx_scan_voutp01,
     oclk_srclkout, oclkb_srclkout, odat_async_fsrdin, osdrin_odat0,
     osdrin_odat1, pcs_clk, pcs_clkb, resetb_sync_buf,
     shift_en_srcclkinn, shift_en_ssrdout, shift_en_ssrldout,
     shift_en_vinp0, shift_en_voutp00, shift_en_voutp01,
     iopad_avmm1_in, iopad_avmm1_out, iopad_clkn, iopad_clkp,
     iopad_inclkn, iopad_inclkp, iopad_sdr_in, iopad_sdr_out,
     avmm1_idat0, avmm1_idat1, avmm1_rstb, avmm_tx_clk_in, clkdr_xr1l,
     clkdr_xr1r, clkdr_xr2l, clkdr_xr2r, clkdr_xr3l, clkdr_xr3r,
     clkdr_xr4l, clkdr_xr4r, iasyncdata_oshared2, idat0_clkn,
     idat0_clkp, idat0_voutp10, idat0_voutp11, idat1_clkn, idat1_clkp,
     idat1_voutp10, idat1_voutp11, idataselb, idataselb_oshared2,
     idataselb_voutp10, idataselb_voutp11, indrv_r12, indrv_r34,
     ipdrv_r12, ipdrv_r34, irxen_inpshared4, irxen_ptxclkin, irxen_r0,
     irxen_r1, irxen_r2, isdrin_idat0, isdrin_idat1, itxen,
     itxen_oshared2, itxen_voutp10, itxen_voutp11,
     jtag_clkdr_in_dirin5, jtag_clkdr_in_voutp10,
     jtag_clkdr_inpshared4, jtag_clkdr_oshared2, jtag_clkdr_ptxclkin,
     jtag_clkdr_ptxclkinn, jtag_clksel, jtag_intest, jtag_mode_in,
     jtag_rstb, jtag_rstb_en, jtag_rx_scan_in_dirin5,
     jtag_rx_scan_in_voutp10, jtag_rx_scan_inpshared4,
     jtag_rx_scan_oshared2, jtag_rx_scan_ptxclkin,
     jtag_rx_scan_ptxclkinn, jtag_tx_scanen_in, jtag_weakpdn,
     jtag_weakpu, oclkn_vinp1, odat0_outpclk1_1, odat1_outpclk1_1,
     rx_shift_en, shift_en_inpshared4, shift_en_oshared2,
     shift_en_ptxclkin, shift_en_ptxclkinn, shift_en_voutp10,
     shift_en_voutp11, vccl_aibnd, vssl_aibnd );

output  avmm1_odat0, avmm1_odat1, avmm2_rx_distclk, avmm2_rx_strbclk,
     avmm2_tx_launch_clk_l0, avmm2_tx_launch_clk_l1, iclkin_dist_vinp0,
     iclkin_dist_vinp1, idat0_voutp00, idat0_voutp01, idat1_voutp00,
     idat1_voutp01, idata0_ssrdout, idata0_ssrldout, idata1_ssrdout,
     idata1_ssrldout, idataselb_ssrdout, idataselb_ssrldout,
     idataselb_voutp00, idataselb_voutp01, ilaunch_clk_ssrdout,
     ilaunch_clk_ssrldout, ilaunch_clk_voutp00, ilaunch_clk_voutp01,
     istrbclk_vinp0, istrbclk_vinp1, itxen_ssrdout, itxen_ssrldout,
     itxen_voutp00, itxen_voutp01, jtag_clkdr_in_srcclkinn,
     jtag_clkdr_in_ssrdout, jtag_clkdr_in_ssrldout, jtag_clkdr_vinp0,
     jtag_clkdr_voutp00, jtag_clkdr_voutp01, jtag_rx_scan_in_srcclkinn,
     jtag_rx_scan_in_ssrdout, jtag_rx_scan_in_ssrldout,
     jtag_rx_scan_vinp0, jtag_rx_scan_voutp00, jtag_rx_scan_voutp01,
     oclk_srclkout, oclkb_srclkout, odat_async_fsrdin, pcs_clk,
     pcs_clkb, resetb_sync_buf, shift_en_srcclkinn, shift_en_ssrdout,
     shift_en_ssrldout, shift_en_vinp0, shift_en_voutp00,
     shift_en_voutp01;

inout  iopad_avmm1_in, iopad_clkn, iopad_clkp, iopad_inclkn,
     iopad_inclkp;

input  avmm1_rstb, avmm_tx_clk_in, clkdr_xr1l, clkdr_xr1r, clkdr_xr2l,
     clkdr_xr2r, clkdr_xr3l, clkdr_xr3r, clkdr_xr4l, clkdr_xr4r,
     iasyncdata_oshared2, idat0_clkn, idat0_clkp, idat0_voutp10,
     idat0_voutp11, idat1_clkn, idat1_clkp, idat1_voutp10,
     idat1_voutp11, idataselb_oshared2, idataselb_voutp10,
     idataselb_voutp11, itxen_oshared2, itxen_voutp10, itxen_voutp11,
     jtag_clkdr_in_dirin5, jtag_clkdr_in_voutp10,
     jtag_clkdr_inpshared4, jtag_clkdr_oshared2, jtag_clkdr_ptxclkin,
     jtag_clkdr_ptxclkinn, jtag_clksel, jtag_intest, jtag_mode_in,
     jtag_rstb, jtag_rstb_en, jtag_rx_scan_in_dirin5,
     jtag_rx_scan_in_voutp10, jtag_rx_scan_inpshared4,
     jtag_rx_scan_oshared2, jtag_rx_scan_ptxclkin,
     jtag_rx_scan_ptxclkinn, jtag_tx_scanen_in, jtag_weakpdn,
     jtag_weakpu, oclkn_vinp1, odat0_outpclk1_1, odat1_outpclk1_1,
     shift_en_inpshared4, shift_en_oshared2, shift_en_ptxclkin,
     shift_en_ptxclkinn, shift_en_voutp10, shift_en_voutp11,
     vccl_aibnd, vssl_aibnd;

output [2:0]  irxen_vinp0;
output [3:0]  osdrin_odat1;
output [3:0]  osdrin_odat0;

inout [1:0]  iopad_avmm1_out;
inout [3:0]  iopad_sdr_in;
inout [3:0]  iopad_sdr_out;

input [1:0]  indrv_r12;
input [1:0]  indrv_r34;
input [1:0]  ipdrv_r34;
input [2:0]  irxen_inpshared4;
input [1:0]  avmm1_idat1;
input [2:0]  itxen;
input [1:0]  avmm1_idat0;
input [2:0]  irxen_ptxclkin;
input [2:0]  irxen_r1;
input [2:0]  irxen_r0;
input [2:0]  idataselb;
input [2:0]  irxen_r2;
input [1:0]  ipdrv_r12;
input [3:0]  isdrin_idat1;
input [3:0]  isdrin_idat0;
input [14:0]  rx_shift_en;

wire clk_distclk_b_nc, clk_distclk, clk_mimic01_b_nc, clk_mimic01, clk_mimic11_b_nc, clk_mimic11, avmm_pcs_clk, avmm_pcs_clk_buf; // Conversion Sript Generated

wire oclk_inclkpb_ext;
// Buses in the design

wire  [0:7]  rx_distclk_l;

wire  [0:7]  rx_distclk_r;

wire  [0:7]  tx_launch_clk_l;

wire  [0:7]  tx_launch_clk_r;


// specify 
//     specparam CDS_LIBNAME  = "aibnd_lib";
//     specparam CDS_CELLNAME = "aibnd_avmm1";
//     specparam CDS_VIEWNAME = "schematic";
// endspecify

aibnd_clktree_avmm  xout_clktree ( /*.vcc_aibnd(vccl_aibnd),
     .vss_aibnd(vssl_aibnd),*/ .lstrbclk_mimic2(nc_clk_mimic),
     .lstrbclk_r_7(tx_launch_clk_r[7]),
     .lstrbclk_r_6(tx_launch_clk_r[6]),
     .lstrbclk_r_5(tx_launch_clk_r[5]),
     .lstrbclk_r_4(tx_launch_clk_r[4]),
     .lstrbclk_r_3(tx_launch_clk_r[3]),
     .lstrbclk_r_2(tx_launch_clk_r[2]),
     .lstrbclk_r_1(tx_launch_clk_r[1]),
     .lstrbclk_r_0(tx_launch_clk_r[0]),
     .lstrbclk_mimic1(nc_clk_mimic1), .lstrbclk_mimic0(nc_clk_mimic0),
     .lstrbclk_l_0(tx_launch_clk_l[0]),
     .lstrbclk_l_1(tx_launch_clk_l[1]),
     .lstrbclk_l_2(tx_launch_clk_l[2]),
     .lstrbclk_l_3(tx_launch_clk_l[3]),
     .lstrbclk_l_4(tx_launch_clk_l[4]),
     .lstrbclk_l_5(tx_launch_clk_l[5]),
     .lstrbclk_l_6(tx_launch_clk_l[6]),
     .lstrbclk_l_7(tx_launch_clk_l[7]), .lstrbclk_rep(nc_clk_rep),
     .clkin(avmm_tx_clk_in_dly));
assign clk_distclk_b_nc = !clk_distclk;

assign clk_mimic01_b_nc = !clk_mimic01;

assign clk_mimic11_b_nc = !clk_mimic11;

aibnd_aliasd  aliasd6 ( .MINUS(ilaunch_clk_voutp01),      .PLUS(tx_launch_clk_l[6]));
aibnd_aliasd  aliasd2 ( .MINUS(idataselb_voutp00), .PLUS(idataselb[0]));
aibnd_aliasd  aliasd7 ( .MINUS(idataselb_voutp01), .PLUS(idataselb[0]));
aibnd_aliasd  aliasv33 ( .MINUS(ilaunch_clk_ssrldout),      .PLUS(tx_launch_clk_r[6]));
aibnd_aliasd  aliasd4 ( .MINUS(itxen_voutp00), .PLUS(itxen[0]));
aibnd_aliasd  aliasd5 ( .MINUS(itxen_voutp01), .PLUS(itxen[0]));
aibnd_aliasd  aliasd15 ( .MINUS(shift_en_ssrdout), .PLUS(rx_shift_en[7]));
aibnd_aliasd  aliasv62 ( .MINUS(iclkin_dist_vinp0), .PLUS(rx_distclk_l[3]));
aibnd_aliasd  aliasv36 ( .MINUS(itxen_ssrldout), .PLUS(itxen[2]));
aibnd_aliasd  aliasv63 ( .MINUS(avmm2_tx_launch_clk_l0),      .PLUS(tx_launch_clk_l[0]));
aibnd_aliasd  aliasv60 ( .MINUS(avmm2_rx_strbclk), .PLUS(rx_distclk_l[6]));
aibnd_aliasd  aliasv61 ( .MINUS(avmm2_rx_distclk), .PLUS(rx_distclk_l[6]));
aibnd_aliasd  aliasv32 ( .MINUS(idataselb_ssrldout), .PLUS(idataselb[2]));
aibnd_aliasd  aliasd11 ( .MINUS(shift_en_srcclkinn), .PLUS(rx_shift_en[4]));
aibnd_aliasd  aliasd14 ( .MINUS(shift_en_ssrldout), .PLUS(rx_shift_en[14]));
aibnd_aliasd  aliasv31 ( .MINUS(ilaunch_clk_ssrdout),      .PLUS(tx_launch_clk_r[7]));
aibnd_aliasd  aliasv0 ( .MINUS(tx_clkn), .PLUS(tx_launch_clk_r[4]));
aibnd_aliasd  aliasv24[2:0] ( .MINUS(irxen_vinp0[2:0]),      .PLUS(irxen_r0[2:0]));
aibnd_aliasd  aliasd13 ( .MINUS(shift_en_voutp01), .PLUS(rx_shift_en[11]));
aibnd_aliasd  aliasd12 ( .MINUS(shift_en_voutp00), .PLUS(rx_shift_en[10]));
aibnd_aliasd  aliasd16 ( .MINUS(istrbclk_vinp1), .PLUS(rx_distclk_l[2]));
aibnd_aliasd  aliasd17 ( .MINUS(iclkin_dist_vinp1), .PLUS(rx_distclk_l[2]));
aibnd_aliasd  aliasv30 ( .MINUS(idataselb_ssrdout), .PLUS(idataselb[2]));
aibnd_aliasd  aliasv64 ( .MINUS(avmm2_tx_launch_clk_l1),      .PLUS(tx_launch_clk_l[1]));
aibnd_aliasd  aliasv25 ( .MINUS(istrbclk_vinp0), .PLUS(rx_distclk_l[3]));
aibnd_aliasd  aliasv1 ( .MINUS(tx_clkp), .PLUS(tx_launch_clk_r[5]));
aibnd_aliasd  aliasd10 ( .MINUS(shift_en_vinp0), .PLUS(rx_shift_en[3]));
aibnd_aliasd  aliasv55 ( .MINUS(itxen_ssrdout), .PLUS(itxen[2]));
aibnd_aliasd  aliasd3 ( .MINUS(ilaunch_clk_voutp00),      .PLUS(tx_launch_clk_l[7]));
aibnd_buffx1_top xtx_clkn ( .idata1_in1_jtag_out(idat1_srcclkoutn),
     .async_dat_in1_jtag_out(nc_async_dat_srcclkoutn),
     .idata0_in1_jtag_out(idat0_srcclkoutn),
     .jtag_clkdr_outn(jtag_clkdr_outn_srcclkoutn),
     .prev_io_shift_en(shift_en_ptxclkinn),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(avmm1_rstb),
     .pd_data_aib(ncdrx_pd_data_out0_txclkn),
     .oclk_out(ncdrx_oclk_txclkp), .oclkb_out(ncdrx_oclkb_txclkp),
     .odat0_out(ncdrx_odat0_txclkp), .odat1_out(ncdrx_odat1_txclkp),
     .odat_async_out(ncdrx_odat_async_txclkp),
     .pd_data_out(ncdrx_pd_data_txclkp), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_srcclkoutn),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0_clkn),
     .idata0_in1(vssl_aibnd), .idata1_in0(idat1_clkn),
     .idata1_in1(vssl_aibnd), .idataselb_in0(idataselb[1]),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(tx_clkn),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r34[1:0]),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0(ipdrv_r34[1:0]),
     .ipdrv_in1({vssl_aibnd, vssl_aibnd}), .irxen_in0({vssl_aibnd,
     vccl_aibnd, vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .istrbclk_in0(jtag_clkdr_outn_srcclkoutn),
     .istrbclk_in1(vssl_aibnd), .itxen_in0(itxen[1]),
     .itxen_in1(vssl_aibnd), .oclk_in1(vssl_aibnd),
     .odat_async_aib(ncdrx_odat_async_out0_txclkn),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[12]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(resetb_sync_buf),
     .jtag_clkdr_out(jtag_clkdr_srcclkoutn),
     .odat1_aib(ncdrx_odat1_out0_txclkn),
     .jtag_rx_scan_out(jtag_rx_scan_srcclkoutn),
     .odat0_aib(ncdrx_odat0_out0_txclkn),
     .oclk_aib(ncdrx_oclk_out0_txclkn),
     .last_bs_out(last_bs_out_dirout3),
     .oclkb_aib(ncdrx_oclkb_out0_txclkn), .jtag_clkdr_in(clkdr_xr4r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_ptxclkinn),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_clkn), .oclkn(oclkn_srcclkoutn), .iclkn(vssl_aibnd),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xavmm1_out1 ( .idata1_in1_jtag_out(idat1_voutp01),
     .async_dat_in1_jtag_out(nc_async_dat_voutp01),
     .idata0_in1_jtag_out(idat0_voutp01),
     .jtag_clkdr_outn(jtag_clkdr_outn_voutp01),
     .prev_io_shift_en(shift_en_voutp11), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(avmm1_rstb), .pd_data_aib(nc_pd_data_avmout01),
     .oclk_out(nc_oclk_avmout1), .oclkb_out(nc_oclkb_avmout1),
     .odat0_out(nc_odat0_avmout1), .odat1_out(nc_odat1_avmout1),
     .odat_async_out(nc_odat_async_avmout1),
     .pd_data_out(nc_pd_data_avmout1), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_voutp01),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(avmm1_idat0[1]),
     .idata0_in1(idat0_voutp11), .idata1_in0(avmm1_idat1[1]),
     .idata1_in1(idat1_voutp11), .idataselb_in0(idataselb[0]),
     .idataselb_in1(idataselb_voutp11), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(tx_launch_clk_l[2]),
     .ilaunch_clk_in1(tx_launch_clk_l[2]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r34[1:0]),
     .indrv_in1(indrv_r34[1:0]), .ipdrv_in0(ipdrv_r34[1:0]),
     .ipdrv_in1(ipdrv_r34[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_voutp01), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[0]), .itxen_in1(itxen_voutp11),
     .oclk_in1(vssl_aibnd), .odat_async_aib(nc_odat_async_avmout01),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[11]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(resetb_sync_buf), .jtag_clkdr_out(jtag_clkdr_voutp01),
     .odat1_aib(nc_odat1_avmout01),
     .jtag_rx_scan_out(jtag_rx_scan_voutp01),
     .odat0_aib(nc_odat0_avmout01), .oclk_aib(nc_oclk_avmout01),
     .last_bs_out(last_bs_out_voutp01), .oclkb_aib(nc_oclkb_avmout01),
     .jtag_clkdr_in(clkdr_xr4l), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_in_dirin5),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_avmm1_out[1]), .oclkn(nc_oclkn_avmout01),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xsdr_in1 ( .idata1_in1_jtag_out(nc_idat1_fsrldin),
     .async_dat_in1_jtag_out(nc_async_dat_fsrldin),
     .idata0_in1_jtag_out(nc_idat0_fsrldin),
     .jtag_clkdr_outn(jtag_clkdr_outn_fsrldin),
     .prev_io_shift_en(shift_en_oshared2), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(avmm1_rstb), .pd_data_aib(nc_pd0_data_fsrldin),
     .oclk_out(nc_oclk_fsrldin), .oclkb_out(nc_oclkb_fsrldin),
     .odat0_out(osdrin_odat0[1]), .odat1_out(osdrin_odat1[1]),
     .odat_async_out(nc_odat_async_fsrldin),
     .pd_data_out(nc_pd_data_fsrldin), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(iasyncdata_oshared2),
     .iclkin_dist_in0(rx_distclk_r[2]), .iclkin_dist_in1(vssl_aibnd),
     .idata0_in0(vssl_aibnd), .idata0_in1(vssl_aibnd),
     .idata1_in0(vssl_aibnd), .idata1_in1(vssl_aibnd),
     .idataselb_in0(vccl_aibnd), .idataselb_in1(idataselb_oshared2),
     .iddren_in0(vssl_aibnd), .iddren_in1(vssl_aibnd),
     .ilaunch_clk_in0(vssl_aibnd), .ilaunch_clk_in1(vssl_aibnd),
     .ilpbk_dat_in0(vssl_aibnd), .ilpbk_dat_in1(vssl_aibnd),
     .ilpbk_en_in0(vssl_aibnd), .ilpbk_en_in1(vssl_aibnd),
     .indrv_in0({vssl_aibnd, vssl_aibnd}), .indrv_in1(indrv_r12[1:0]),
     .ipdrv_in0({vssl_aibnd, vssl_aibnd}), .ipdrv_in1(ipdrv_r12[1:0]),
     .irxen_in0(irxen_r2[2:0]), .irxen_in1({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .istrbclk_in0(rx_distclk_r[2]),
     .istrbclk_in1(vssl_aibnd), .itxen_in0(vssl_aibnd),
     .itxen_in1(itxen_oshared2), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_out0_fsrldin),
     .oclkb_in1(vssl_aibnd), .odat0_in1(ossrldin_odat0),
     .odat1_in1(ossrldin_odat1), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[6]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(resetb_sync_buf),
     .jtag_clkdr_out(jtag_clkdr_out_fsrldin),
     .odat1_aib(nc_odat0_out1_fsrldin),
     .jtag_rx_scan_out(jtag_rx_scan_out_fsrldin),
     .odat0_aib(nc_odat0_out0_fsrldin),
     .oclk_aib(nc_oclk_out0_fsrldin),
     .last_bs_out(last_bs_out_fsrldin),
     .oclkb_aib(nc_oclkb_out0_fsrldin), .jtag_clkdr_in(clkdr_xr2r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_oshared2),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_sdr_in[1]), .oclkn(nc_oclkn_out0_fsrldin),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xsdr_in0 ( .idata1_in1_jtag_out(nc_idat1_ssrldin),
     .async_dat_in1_jtag_out(nc_async_dat_ssrldin),
     .idata0_in1_jtag_out(nc_idat0_ssrldin),
     .jtag_clkdr_outn(jtag_clkdr_outn_ssrldin),
     .prev_io_shift_en(rx_shift_en[6]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(avmm1_rstb), .pd_data_aib(nc_pd_data_out0_ssrldin),
     .oclk_out(nc_oclk_ssrldin), .oclkb_out(nc_oclkb_ssrldin),
     .odat0_out(osdrin_odat0[0]), .odat1_out(osdrin_odat1[0]),
     .odat_async_out(nc_odat_async_ssrldin),
     .pd_data_out(nc_pd_data_ssrldin), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_r[0]),
     .iclkin_dist_in1(rx_distclk_r[2]), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r2[2:0]), .irxen_in1(irxen_r2[2:0]),
     .istrbclk_in0(rx_distclk_r[0]), .istrbclk_in1(rx_distclk_r[0]),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_out0_ssrldin),
     .oclkb_in1(vssl_aibnd), .odat0_in1(odat0_srcclkinn),
     .odat1_in1(odat1_srcclkinn), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[5]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(resetb_sync_buf),
     .jtag_clkdr_out(jtag_clkdr_out_ssrldin),
     .odat1_aib(ossrldin_odat1),
     .jtag_rx_scan_out(jtag_rx_scan_out_ssrldin),
     .odat0_aib(ossrldin_odat0), .oclk_aib(nc_oclk_out0_ssrldin),
     .last_bs_out(last_bs_out_ssrldin),
     .oclkb_aib(nc_oclkb_out0_ssrldin), .jtag_clkdr_in(clkdr_xr2r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_fsrldin),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_sdr_in[0]), .oclkn(nc_oclkn_out0_ssrldin),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xrx_clkn ( .idata1_in1_jtag_out(nc_idat1_srcclkinn),
     .async_dat_in1_jtag_out(nc_async_dat_srcclkinn),
     .idata0_in1_jtag_out(nc_idat0_srcclkinn),
     .jtag_clkdr_outn(jtag_clkdr_outn_srcclkinn),
     .prev_io_shift_en(rx_shift_en[5]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(avmm1_rstb), .pd_data_aib(pd_data_srcclkinn),
     .oclk_out(oclk_inclkn), .oclkb_out(oclk_inclknb),
     .odat0_out(ncdrx_odat0_inclkn), .odat1_out(ncdrx_odat1_inclkn),
     .odat_async_out(odirectin_data_inclkn),
     .pd_data_out(pd_data_inclkn), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_r[4]),
     .iclkin_dist_in1(rx_distclk_r[0]), .idata0_in0(vccl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .irxen_in1(irxen_r2[2:0]), .istrbclk_in0(rx_distclk_r[4]),
     .istrbclk_in1(rx_distclk_r[4]), .itxen_in0(vssl_aibnd),
     .itxen_in1(vssl_aibnd), .oclk_in1(vssl_aibnd),
     .odat_async_aib(odirectin_data_srcclkinn), .oclkb_in1(vssl_aibnd),
     .odat0_in1(vssl_aibnd), .odat1_in1(vssl_aibnd),
     .odat_async_in1(vssl_aibnd), .shift_en(rx_shift_en[4]),
     .pd_data_in1(vssl_aibnd), .dig_rstb(resetb_sync_buf),
     .jtag_clkdr_out(jtag_clkdr_in_srcclkinn),
     .odat1_aib(odat1_srcclkinn),
     .jtag_rx_scan_out(jtag_rx_scan_in_srcclkinn),
     .odat0_aib(odat0_srcclkinn), .oclk_aib(nc_oclk_srcclkinn),
     .last_bs_out(nc), .oclkb_aib(nc_oclkb_srcclkinn),
     .jtag_clkdr_in(clkdr_xr2r), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_out_ssrldin),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_inclkn), .oclkn(oclkn_inclkn), .iclkn(vssl_aibnd),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xtx_clkp ( .idata1_in1_jtag_out(idat1_srclkout),
     .async_dat_in1_jtag_out(nc_async_dat_srclkout),
     .idata0_in1_jtag_out(idat0_srclkout),
     .jtag_clkdr_outn(jtag_clkdr_outn_srclkout),
     .prev_io_shift_en(shift_en_ptxclkin), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(avmm1_rstb), .pd_data_aib(ncdrx_pd_data_out0_txclkp),
     .oclk_out(ncdrx_oclk_txclkp1), .oclkb_out(ncdrx_oclkb_txclkp1),
     .odat0_out(ncdrx_odat0_txclkp1), .odat1_out(ncdrx_odat1_txclkp1),
     .odat_async_out(ncdrx_odat_async_txclkp1),
     .pd_data_out(ncdrx_pd_data_txclkp1), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_srclkout),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(idat0_clkp),
     .idata0_in1(vssl_aibnd), .idata1_in0(idat1_clkp),
     .idata1_in1(vssl_aibnd), .idataselb_in0(idataselb[1]),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(tx_clkp),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r34[1:0]),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0(ipdrv_r34[1:0]),
     .ipdrv_in1({vssl_aibnd, vssl_aibnd}), .irxen_in0({vssl_aibnd,
     vccl_aibnd, vssl_aibnd}), .irxen_in1(irxen_ptxclkin[2:0]),
     .istrbclk_in0(jtag_clkdr_outn_srclkout),
     .istrbclk_in1(vssl_aibnd), .itxen_in0(itxen[1]),
     .itxen_in1(vssl_aibnd), .oclk_in1(vssl_aibnd),
     .odat_async_aib(ncdrx_odat_async_out0_txclkp),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[9]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(resetb_sync_buf), .jtag_clkdr_out(jtag_clkdr_srclkout),
     .odat1_aib(ncdrx_odat1_out0_txclkp),
     .jtag_rx_scan_out(jtag_rx_scan_srclkout),
     .odat0_aib(ncdrx_odat0_out0_txclkp), .oclk_aib(oclk_srclkout),
     .last_bs_out(last_bs_out_directout0), .oclkb_aib(oclkb_srclkout),
     .jtag_clkdr_in(clkdr_xr3r), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_ptxclkin),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_clkp), .oclkn(ncdrx_oclkn_txclkp),
     .iclkn(oclkn_srcclkoutn), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xsdr_out1 ( .idata1_in1_jtag_out(idat1_fsrdout),
     .async_dat_in1_jtag_out(nc_async_dat_fsrdout),
     .idata0_in1_jtag_out(idat0_fsrdout),
     .jtag_clkdr_outn(jtag_clkdr_outn_fsrdout),
     .prev_io_shift_en(rx_shift_en[12]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(avmm1_rstb), .pd_data_aib(nc_pd_data_out0_fsrlout),
     .oclk_out(nc_oclk_fsrout), .oclkb_out(nc_oclkb_fsrout),
     .odat0_out(nc_odat0_fsrout), .odat1_out(nc_odat1_fsrout),
     .odat_async_out(nc_odat_async_fsrout),
     .pd_data_out(nc_pd_data_fsrout), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_fsrdout),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(isdrin_idat0[1]),
     .idata0_in1(idat0_srcclkoutn), .idata1_in0(isdrin_idat1[1]),
     .idata1_in1(idat1_srcclkoutn), .idataselb_in0(idataselb[2]),
     .idataselb_in1(idataselb[1]), .iddren_in0(vssl_aibnd),
     .iddren_in1(vccl_aibnd), .ilaunch_clk_in0(tx_launch_clk_r[0]),
     .ilaunch_clk_in1(tx_launch_clk_r[0]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r34[1:0]),
     .indrv_in1(indrv_r34[1:0]), .ipdrv_in0(ipdrv_r34[1:0]),
     .ipdrv_in1(ipdrv_r34[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_fsrdout), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[2]), .itxen_in1(itxen[1]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_out0_fsrlout),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[13]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(resetb_sync_buf),
     .jtag_clkdr_out(jtag_clkdr_out_fsrdout),
     .odat1_aib(nc_odat1_out0_fsrlout),
     .jtag_rx_scan_out(jtag_rx_scan_out_fsrdout),
     .odat0_aib(nc_odat0_out0_fsrlout),
     .oclk_aib(nc_oclk_out0_fsrlout),
     .last_bs_out(last_bs_out_fsrdout),
     .oclkb_aib(nc_oclkb_out0_fsrlout), .jtag_clkdr_in(clkdr_xr4r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_srcclkoutn),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_sdr_out[1]), .oclkn(nc_oclkn_out0_fsrlout),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xsdr_out0 ( .idata1_in1_jtag_out(idata1_ssrldout),
     .async_dat_in1_jtag_out(nc_async_dat_ssrldout),
     .idata0_in1_jtag_out(idata0_ssrldout),
     .jtag_clkdr_outn(jtag_clkdr_outn_ssrldout),
     .prev_io_shift_en(rx_shift_en[13]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(avmm1_rstb), .pd_data_aib(nc_pd_data_out0_ssrldrout),
     .oclk_out(nc_oclk_ssrldout), .oclkb_out(nc_oclkb_ssrldout),
     .odat0_out(nc_odat0_ssrldout), .odat1_out(nc_odat1_ssrldout),
     .odat_async_out(nc_odat_async_ssrldout),
     .pd_data_out(nc_pd_data_ssrldout), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_ssrldout),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(isdrin_idat0[0]),
     .idata0_in1(idat0_fsrdout), .idata1_in0(isdrin_idat1[0]),
     .idata1_in1(idat1_fsrdout), .idataselb_in0(idataselb[2]),
     .idataselb_in1(idataselb[2]), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(tx_launch_clk_r[2]),
     .ilaunch_clk_in1(tx_launch_clk_r[2]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r34[1:0]),
     .indrv_in1(indrv_r34[1:0]), .ipdrv_in0(ipdrv_r34[1:0]),
     .ipdrv_in1(ipdrv_r34[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_ssrldout),
     .istrbclk_in1(vssl_aibnd), .itxen_in0(itxen[2]),
     .itxen_in1(itxen[2]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_out0_ssrldrout),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[14]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(resetb_sync_buf),
     .jtag_clkdr_out(jtag_clkdr_in_ssrldout),
     .odat1_aib(nc_odat1_out0_ssrldrout),
     .jtag_rx_scan_out(jtag_rx_scan_in_ssrldout),
     .odat0_aib(nc_odat0_out0_ssrldrout),
     .oclk_aib(nc_oclk_out0_ssrldrout),
     .last_bs_out(last_bs_out_ssrldout),
     .oclkb_aib(nc_oclkb_out0_ssrldrout), .jtag_clkdr_in(clkdr_xr4r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_fsrdout),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_out_fsrdout), .iopad(iopad_sdr_out[0]),
     .oclkn(nc_oclkn_out0_ssrldrout), .iclkn(vssl_aibnd),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xsdr_in3 ( .idata1_in1_jtag_out(nc_idat1_fsrdin),
     .async_dat_in1_jtag_out(nc_async_dat_fsrdin),
     .idata0_in1_jtag_out(nc_idat0_fsrdin),
     .jtag_clkdr_outn(jtag_clkdr_outn_fsrdin),
     .prev_io_shift_en(shift_en_inpshared4),
     .jtag_rstb_en(jtag_rstb_en), .jtag_clksel(jtag_clksel),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd),
     .jtag_intest(jtag_intest), .anlg_rstb(avmm1_rstb),
     .pd_data_aib(nc_pd_data_out0_fsrdin), .oclk_out(nc_oclk_fsrdin),
     .oclkb_out(nc_oclkb_fsrdin), .odat0_out(osdrin_odat0[3]),
     .odat1_out(osdrin_odat1[3]),
     .odat_async_out(nc_odat_async_fsrdin),
     .pd_data_out(nc_pd_data_fsrdin), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_r[3]),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r2[2:0]), .irxen_in1(irxen_inpshared4[2:0]),
     .istrbclk_in0(rx_distclk_r[3]), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(odat_async_fsrdin),
     .oclkb_in1(vssl_aibnd), .odat0_in1(ossrdin_odat0),
     .odat1_in1(ossrdin_odat1), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[0]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(resetb_sync_buf),
     .jtag_clkdr_out(jtag_clkdr_out_fsrdin),
     .odat1_aib(nc_odat1_out0_fsrdin),
     .jtag_rx_scan_out(jtag_rx_scan_out_fsrdin),
     .odat0_aib(nc_odat0_out0_fsrdin), .oclk_aib(nc_oclk_out0_fsrdin),
     .last_bs_out(last_bs_out_fsrdin),
     .oclkb_aib(nc_oclkb_out0_fsrdin), .jtag_clkdr_in(clkdr_xr1r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_inpshared4),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_sdr_in[3]), .oclkn(nc_oclkn_out0_fsrdin),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xrx_clkp ( .idata1_in1_jtag_out(nc_idat1_srcclkin),
     .async_dat_in1_jtag_out(nc_async_dat_srcclkin),
     .idata0_in1_jtag_out(nc_idat0_srcclkin),
     .jtag_clkdr_outn(jtag_clkdr_outn_srcclkin),
     .prev_io_shift_en(rx_shift_en[1]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(avmm1_rstb), .pd_data_aib(pd_data_srcclkin),
     .oclk_out(oclk_inclkp), .oclkb_out(oclk_inclkpb),
     .odat0_out(ncdrx_odat0_inclkp), .odat1_out(ncdrx_odat1_inclkp),
     .odat_async_out(odirectin_data_inclkp),
     .pd_data_out(pd_data_inclkp), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_r[5]),
     .iclkin_dist_in1(rx_distclk_r[1]), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vccl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vccl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r1[2:0]), .irxen_in1(irxen_r2[2:0]),
     .istrbclk_in0(rx_distclk_r[5]), .istrbclk_in1(rx_distclk_r[5]),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(oclk_vinp0), .odat_async_aib(odirectin_data_srcclkin),
     .oclkb_in1(oclk_inclkpb_ext), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[2]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(resetb_sync_buf),
     .jtag_clkdr_out(jtag_clkdr_in_srcclkin),
     .odat1_aib(odat1_srcclkin),
     .jtag_rx_scan_out(jtag_rx_scan_in_srcclkin),
     .odat0_aib(odat0_srcclkin), .oclk_aib(ncdrx_oclk_srcclkin),
     .last_bs_out(last_bs_out_srcclkin),
     .oclkb_aib(drx_oclkb_srcclkin), .jtag_clkdr_in(clkdr_xr1r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_ssrdin),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_inclkp), .oclkn(ncdrx_oclkn_srcclkin),
     .iclkn(oclkn_inclkn), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xavmm1_out0 ( .idata1_in1_jtag_out(idat1_voutp00),
     .async_dat_in1_jtag_out(nc_async_dat_voutp00),
     .idata0_in1_jtag_out(idat0_voutp00),
     .jtag_clkdr_outn(jtag_clkdr_outn_voutp00),
     .prev_io_shift_en(shift_en_voutp10), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(avmm1_rstb), .pd_data_aib(nc_pd_data_avmout0),
     .oclk_out(nc_oclk_avmout011), .oclkb_out(nc_oclkb_avmout011),
     .odat0_out(nc_odat0_avmout011), .odat1_out(nc_odat1_avmout011),
     .odat_async_out(nc_odat_async_avmout011),
     .pd_data_out(nc_pd_data_avmout011), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_voutp00),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(avmm1_idat0[0]),
     .idata0_in1(idat0_voutp10), .idata1_in0(avmm1_idat1[0]),
     .idata1_in1(idat1_voutp10), .idataselb_in0(idataselb[0]),
     .idataselb_in1(idataselb_voutp10), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(tx_launch_clk_l[3]),
     .ilaunch_clk_in1(tx_launch_clk_l[3]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r34[1:0]),
     .indrv_in1(indrv_r34[1:0]), .ipdrv_in0(ipdrv_r34[1:0]),
     .ipdrv_in1(ipdrv_r34[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_voutp00), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[0]), .itxen_in1(itxen_voutp10),
     .oclk_in1(vssl_aibnd), .odat_async_aib(nc_odat_async_avmout0),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[10]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(resetb_sync_buf), .jtag_clkdr_out(jtag_clkdr_voutp00),
     .odat1_aib(nc_odat1_avmout0),
     .jtag_rx_scan_out(jtag_rx_scan_voutp00),
     .odat0_aib(nc_odat0_avmout0), .oclk_aib(nc_oclk_avmout0),
     .last_bs_out(last_bs_out_voutp00), .oclkb_aib(nc_oclkb_avmout0),
     .jtag_clkdr_in(clkdr_xr3l), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_in_voutp10),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_avmm1_out[0]), .oclkn(nc_oclkn_avmout0),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xsdr_out3 ( .idata1_in1_jtag_out(idat1_fsrldout),
     .async_dat_in1_jtag_out(nc_async_dat_fsrldout),
     .idata0_in1_jtag_out(idat0_fsrldout),
     .jtag_clkdr_outn(jtag_clkdr_outn_fsrldout),
     .prev_io_shift_en(rx_shift_en[9]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(avmm1_rstb), .pd_data_aib(nc_pd_data_out0_fsrout),
     .oclk_out(nc_oclk_fsrout1), .oclkb_out(nc_oclkb_fsrout1),
     .odat0_out(nc_odat0_fsrout1), .odat1_out(nc_odat1_fsrout1),
     .odat_async_out(nc_odat_async_fsrout1),
     .pd_data_out(nc_pd_data_fsrout1), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_fsrldout),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(isdrin_idat0[3]),
     .idata0_in1(idat0_srclkout), .idata1_in0(isdrin_idat1[3]),
     .idata1_in1(idat1_srclkout), .idataselb_in0(idataselb[2]),
     .idataselb_in1(idataselb[1]), .iddren_in0(vssl_aibnd),
     .iddren_in1(vccl_aibnd), .ilaunch_clk_in0(tx_launch_clk_r[1]),
     .ilaunch_clk_in1(tx_launch_clk_r[1]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r34[1:0]),
     .indrv_in1(indrv_r34[1:0]), .ipdrv_in0(ipdrv_r34[1:0]),
     .ipdrv_in1(ipdrv_r34[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_fsrldout),
     .istrbclk_in1(vssl_aibnd), .itxen_in0(itxen[2]),
     .itxen_in1(itxen[1]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_out0_fsrout),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[8]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(resetb_sync_buf),
     .jtag_clkdr_out(jtag_clkdr_out_fsrldout),
     .odat1_aib(nc_odat1_out0_fsrout),
     .jtag_rx_scan_out(jtag_rx_scan_out_fsrldout),
     .odat0_aib(nc_odat0_out0_fsrout), .oclk_aib(nc_oclk_out0_fsrout),
     .last_bs_out(last_bs_out_fsrldout),
     .oclkb_aib(nc_oclkb_out0_fsrout), .jtag_clkdr_in(clkdr_xr3r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_srclkout),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_sdr_out[3]), .oclkn(nc_oclkn_out0_fsrout),
     .iclkn(vssl_aibnd), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xsdr_in2 ( .idata1_in1_jtag_out(nc_idat1_ssrdin),
     .async_dat_in1_jtag_out(nc_async_dat_ssrdin),
     .idata0_in1_jtag_out(nc_idat0_ssrdin),
     .jtag_clkdr_outn(jtag_clkdr_outn_ssrdin),
     .prev_io_shift_en(rx_shift_en[0]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(avmm1_rstb), .pd_data_aib(nc_pd_data_out0_ssrdin),
     .oclk_out(nc_oclk_ssrdin), .oclkb_out(nc_oclkb_ssrdin),
     .odat0_out(osdrin_odat0[2]), .odat1_out(osdrin_odat1[2]),
     .odat_async_out(nc_odat_async_ssrdin),
     .pd_data_out(nc_pd_data_ssrdin), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd), .iclkin_dist_in0(rx_distclk_r[1]),
     .iclkin_dist_in1(rx_distclk_r[3]), .idata0_in0(vssl_aibnd),
     .idata0_in1(vssl_aibnd), .idata1_in0(vssl_aibnd),
     .idata1_in1(vssl_aibnd), .idataselb_in0(vccl_aibnd),
     .idataselb_in1(vssl_aibnd), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(vssl_aibnd),
     .ilaunch_clk_in1(vssl_aibnd), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0({vssl_aibnd, vssl_aibnd}),
     .indrv_in1({vssl_aibnd, vssl_aibnd}), .ipdrv_in0({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in1({vssl_aibnd, vssl_aibnd}),
     .irxen_in0(irxen_r2[2:0]), .irxen_in1(irxen_r2[2:0]),
     .istrbclk_in0(rx_distclk_r[1]), .istrbclk_in1(rx_distclk_r[1]),
     .itxen_in0(vssl_aibnd), .itxen_in1(vssl_aibnd),
     .oclk_in1(vssl_aibnd), .odat_async_aib(nc_odat_async_out0_ssrdin),
     .oclkb_in1(vssl_aibnd), .odat0_in1(odat0_srcclkin),
     .odat1_in1(odat1_srcclkin), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[1]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(resetb_sync_buf),
     .jtag_clkdr_out(jtag_clkdr_out_ssrdin), .odat1_aib(ossrdin_odat1),
     .jtag_rx_scan_out(jtag_rx_scan_out_ssrdin),
     .odat0_aib(ossrdin_odat0), .oclk_aib(nc_oclk_out0_ssrdin),
     .last_bs_out(last_bs_out_ssrdin),
     .oclkb_aib(nc_oclkb_out0_ssrdin), .jtag_clkdr_in(clkdr_xr1r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_fsrdin),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_sdr_in[2]), .oclkn(nc_oclkn_out0_ssrdin),
     .test_weakpd(jtag_weakpdn), .iclkn(vssl_aibnd),
     .test_weakpu(jtag_weakpu));
aibnd_buffx1_top xrx ( .idata1_in1_jtag_out(nc_idat1_vinp0),
     .async_dat_in1_jtag_out(nc_async_dat_vinp0),
     .idata0_in1_jtag_out(nc_idat0_vinp0),
     .jtag_clkdr_outn(jtag_clkdr_outn_vinp0),
     .prev_io_shift_en(rx_shift_en[2]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(avmm1_rstb), .pd_data_aib(nc_pd_data_out0_rx),
     .oclk_out(nc_oclk_rx), .oclkb_out(nc_oclkb_rx),
     .odat0_out(avmm1_odat0), .odat1_out(avmm1_odat1),
     .odat_async_out(nc_odat_async_rx), .pd_data_out(nc_pd_data_rx),
     .async_dat_in0(vssl_aibnd), .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(rx_distclk_l[7]), .iclkin_dist_in1(vssl_aibnd),
     .idata0_in0(vssl_aibnd), .idata0_in1(vssl_aibnd),
     .idata1_in0(vssl_aibnd), .idata1_in1(vssl_aibnd),
     .idataselb_in0(vccl_aibnd), .idataselb_in1(vssl_aibnd),
     .iddren_in0(vssl_aibnd), .iddren_in1(vssl_aibnd),
     .ilaunch_clk_in0(vssl_aibnd), .ilaunch_clk_in1(vssl_aibnd),
     .ilpbk_dat_in0(vssl_aibnd), .ilpbk_dat_in1(vssl_aibnd),
     .ilpbk_en_in0(vssl_aibnd), .ilpbk_en_in1(vssl_aibnd),
     .indrv_in0({vssl_aibnd, vssl_aibnd}), .indrv_in1({vssl_aibnd,
     vssl_aibnd}), .ipdrv_in0({vssl_aibnd, vssl_aibnd}),
     .ipdrv_in1({vssl_aibnd, vssl_aibnd}), .irxen_in0(irxen_r0[2:0]),
     .irxen_in1(irxen_r1[2:0]), .istrbclk_in0(rx_distclk_l[7]),
     .istrbclk_in1(vssl_aibnd), .itxen_in0(vssl_aibnd),
     .itxen_in1(vssl_aibnd), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_out0_rx), .oclkb_in1(vssl_aibnd),
     .odat0_in1(odat0_outpclk1_1), .odat1_in1(odat1_outpclk1_1),
     .odat_async_in1(vssl_aibnd), .shift_en(rx_shift_en[3]),
     .pd_data_in1(vssl_aibnd), .dig_rstb(resetb_sync_buf),
     .jtag_clkdr_out(jtag_clkdr_vinp0), .odat1_aib(nc_odat1_out0_rx),
     .jtag_rx_scan_out(jtag_rx_scan_vinp0),
     .odat0_aib(nc_odat0_out0_rx), .oclk_aib(oclk_vinp0),
     .last_bs_out(last_bs_out_vinp0), .oclkb_aib(oclkb_vinp0),
     .jtag_clkdr_in(clkdr_xr1l), .jtag_mode_in(jtag_mode_in),
     .jtag_rstb(jtag_rstb), .jtag_tx_scan_in(jtag_rx_scan_in_srcclkin),
     .jtag_tx_scanen_in(jtag_tx_scanen_in), .last_bs_in(vssl_aibnd),
     .iopad(iopad_avmm1_in), .oclkn(nc_oclkn_out0_rx),
     .iclkn(oclkn_vinp1), .test_weakpu(jtag_weakpu),
     .test_weakpd(jtag_weakpdn));
aibnd_buffx1_top xsdr_out2 ( .idata1_in1_jtag_out(idata1_ssrdout),
     .async_dat_in1_jtag_out(nc_async_dat_ssrdout),
     .idata0_in1_jtag_out(idata0_ssrdout),
     .jtag_clkdr_outn(jtag_clkdr_outn_ssrdout),
     .prev_io_shift_en(rx_shift_en[8]), .jtag_rstb_en(jtag_rstb_en),
     .jtag_clksel(jtag_clksel), .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .jtag_intest(jtag_intest),
     .anlg_rstb(avmm1_rstb), .pd_data_aib(nc_pd_data_out0_sdrout),
     .oclk_out(nc_oclk_sdrout), .oclkb_out(nc_oclkb_ssdrout),
     .odat0_out(nc_odat0_sdrout), .odat1_out(nc_odat1_ssdrout),
     .odat_async_out(nc_odat_async_sdrout),
     .pd_data_out(nc_pd_data_sdrout), .async_dat_in0(vssl_aibnd),
     .async_dat_in1(vssl_aibnd),
     .iclkin_dist_in0(jtag_clkdr_outn_ssrdout),
     .iclkin_dist_in1(vssl_aibnd), .idata0_in0(isdrin_idat0[2]),
     .idata0_in1(idat0_fsrldout), .idata1_in0(isdrin_idat1[2]),
     .idata1_in1(idat1_fsrldout), .idataselb_in0(idataselb[2]),
     .idataselb_in1(idataselb[2]), .iddren_in0(vssl_aibnd),
     .iddren_in1(vssl_aibnd), .ilaunch_clk_in0(tx_launch_clk_r[3]),
     .ilaunch_clk_in1(tx_launch_clk_r[3]), .ilpbk_dat_in0(vssl_aibnd),
     .ilpbk_dat_in1(vssl_aibnd), .ilpbk_en_in0(vssl_aibnd),
     .ilpbk_en_in1(vssl_aibnd), .indrv_in0(indrv_r34[1:0]),
     .indrv_in1(indrv_r34[1:0]), .ipdrv_in0(ipdrv_r34[1:0]),
     .ipdrv_in1(ipdrv_r34[1:0]), .irxen_in0({vssl_aibnd, vccl_aibnd,
     vssl_aibnd}), .irxen_in1({vssl_aibnd, vccl_aibnd, vssl_aibnd}),
     .istrbclk_in0(jtag_clkdr_outn_ssrdout), .istrbclk_in1(vssl_aibnd),
     .itxen_in0(itxen[2]), .itxen_in1(itxen[2]), .oclk_in1(vssl_aibnd),
     .odat_async_aib(nc_odat_async_out0_sdrout),
     .oclkb_in1(vssl_aibnd), .odat0_in1(vssl_aibnd),
     .odat1_in1(vssl_aibnd), .odat_async_in1(vssl_aibnd),
     .shift_en(rx_shift_en[7]), .pd_data_in1(vssl_aibnd),
     .dig_rstb(resetb_sync_buf),
     .jtag_clkdr_out(jtag_clkdr_in_ssrdout),
     .odat1_aib(nc_odat1_out0_ssdrout),
     .jtag_rx_scan_out(jtag_rx_scan_in_ssrdout),
     .odat0_aib(nc_odat0_out0_sdrout), .oclk_aib(nc_oclk_out0_sdrout),
     .last_bs_out(last_bs_out_ssrdout),
     .oclkb_aib(nc_oclkb_out0_ssdrout), .jtag_clkdr_in(clkdr_xr3r),
     .jtag_mode_in(jtag_mode_in), .jtag_rstb(jtag_rstb),
     .jtag_tx_scan_in(jtag_rx_scan_out_fsrldout),
     .jtag_tx_scanen_in(jtag_tx_scanen_in),
     .last_bs_in(last_bs_out_fsrldout), .iopad(iopad_sdr_out[2]),
     .oclkn(nc_oclkn_out0_ssdrout), .iclkn(vssl_aibnd),
     .test_weakpu(jtag_weakpu), .test_weakpd(jtag_weakpdn));
aibnd_clktree_avmm_pcs  xin_clktree ( /*.vcc_aibnd(vccl_aibnd),
     .vss_aibnd(vssl_aibnd),*/ .lstrbclk_mimic2(clk_distclk),
     .lstrbclk_r_7(rx_distclk_r[7]), .lstrbclk_r_6(rx_distclk_r[6]),
     .lstrbclk_r_5(rx_distclk_r[5]), .lstrbclk_r_4(rx_distclk_r[4]),
     .lstrbclk_r_3(rx_distclk_r[3]), .lstrbclk_r_2(rx_distclk_r[2]),
     .lstrbclk_r_1(rx_distclk_r[1]), .lstrbclk_r_0(rx_distclk_r[0]),
     .lstrbclk_mimic1(clk_mimic11), .lstrbclk_mimic0(clk_mimic01),
     .lstrbclk_l_0(rx_distclk_l[0]), .lstrbclk_l_1(rx_distclk_l[1]),
     .lstrbclk_l_2(rx_distclk_l[2]), .lstrbclk_l_3(rx_distclk_l[3]),
     .lstrbclk_l_4(rx_distclk_l[4]), .lstrbclk_l_5(rx_distclk_l[5]),
     .lstrbclk_l_6(rx_distclk_l[6]), .lstrbclk_l_7(rx_distclk_l[7]),
     .lstrbclk_rep(avmm_pcs_clk), .clkin(oclk_inclkpb_ext));
aibnd_txdat_mimic x570 ( .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .idata_out(avmm_tx_clk_in_dly),
     .idata_in(avmm_tx_clk_in));
assign avmm_pcs_clk_buf = avmm_pcs_clk ;
aibnd_rxdat_mimic x571 ( .odat_out(pcs_clk), .odat_in(pre_pcs_clk),
     .vssl_aibnd(vssl_aibnd), .vccl_aibnd(vccl_aibnd));
aibnd_avmm_rst_sync x568 ( .vssl_aibnd(vssl_aibnd),
     .vccl_aibnd(vccl_aibnd), .pcs_clk(pre_pcs_clk),
     .pcs_clkb(pcs_clkb), .resetb_sync_buf(resetb_sync_buf),
     .avmm_clk(avmm_pcs_clk_buf), .avmm_rstb(avmm1_rstb));


aibnd_clkmux2 xavmm_rx_clkmx ( 
      .oclk_out(oclk_inclkpb_ext),
     .mux_sel(rx_shift_en[2]), .oclk_in0(drx_oclkb_srcclkin),
     .oclk_in1(oclkb_vinp0));

endmodule

