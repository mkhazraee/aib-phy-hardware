// SPDX-License-Identifier: Apache-2.0
// Copyright (C) 2019 Intel Corporation. 
// *****************************************************************************
// *****************************************************************************
//  Copyright © 2016 Altera Corporation.  
// *****************************************************************************
//  Module Name :  c3lib_ecc_dec_c39_d32
//  Date        :  Thu Jan 26 18:03:00 2017
//  Description :  ECC checker (based on the standard Extended Hamming Code
//                 scheme). Code generated by ecc_chk.pl script (command line
//                 options used: -num_data_bits 32).
// *****************************************************************************

module c3lib_ecc_dec_c39_d32(

  output logic		o_int_sec,
  output logic		o_int_ded,
  output logic[ 5 : 0 ]	o_syndrome,

  input  logic[ 38 : 0 ]	i_code,
  output logic[ 31 : 0 ]	o_data

);

// Declarations
logic		parity0;
logic[ 38 : 1 ]	correct_bit;

// Validate parity bits
assign parity0 = i_code[ 0 ] ^ i_code[ 1 ] ^ i_code[ 2 ] ^ i_code[ 3 ] ^ i_code[ 4 ] ^ i_code[ 5 ] ^ i_code[ 6 ] ^ i_code[ 7 ] ^ i_code[ 8 ] ^ i_code[ 9 ] ^ i_code[ 10 ] ^ i_code[ 11 ] ^ i_code[ 12 ] ^ i_code[ 13 ] ^ i_code[ 14 ] ^ i_code[ 15 ] ^ i_code[ 16 ] ^ i_code[ 17 ] ^ i_code[ 18 ] ^ i_code[ 19 ] ^ i_code[ 20 ] ^ i_code[ 21 ] ^ i_code[ 22 ] ^ i_code[ 23 ] ^ i_code[ 24 ] ^ i_code[ 25 ] ^ i_code[ 26 ] ^ i_code[ 27 ] ^ i_code[ 28 ] ^ i_code[ 29 ] ^ i_code[ 30 ] ^ i_code[ 31 ] ^ i_code[ 32 ] ^ i_code[ 33 ] ^ i_code[ 34 ] ^ i_code[ 35 ] ^ i_code[ 36 ] ^ i_code[ 37 ] ^ i_code[ 38 ];
assign o_syndrome[ 0 ] = i_code[ 1 ] ^ i_code[ 3 ] ^ i_code[ 5 ] ^ i_code[ 7 ] ^ i_code[ 9 ] ^ i_code[ 11 ] ^ i_code[ 13 ] ^ i_code[ 15 ] ^ i_code[ 17 ] ^ i_code[ 19 ] ^ i_code[ 21 ] ^ i_code[ 23 ] ^ i_code[ 25 ] ^ i_code[ 27 ] ^ i_code[ 29 ] ^ i_code[ 31 ] ^ i_code[ 33 ] ^ i_code[ 35 ] ^ i_code[ 37 ];
assign o_syndrome[ 1 ] = i_code[ 2 ] ^ i_code[ 3 ] ^ i_code[ 6 ] ^ i_code[ 7 ] ^ i_code[ 10 ] ^ i_code[ 11 ] ^ i_code[ 14 ] ^ i_code[ 15 ] ^ i_code[ 18 ] ^ i_code[ 19 ] ^ i_code[ 22 ] ^ i_code[ 23 ] ^ i_code[ 26 ] ^ i_code[ 27 ] ^ i_code[ 30 ] ^ i_code[ 31 ] ^ i_code[ 34 ] ^ i_code[ 35 ] ^ i_code[ 38 ];
assign o_syndrome[ 2 ] = i_code[ 4 ] ^ i_code[ 5 ] ^ i_code[ 6 ] ^ i_code[ 7 ] ^ i_code[ 12 ] ^ i_code[ 13 ] ^ i_code[ 14 ] ^ i_code[ 15 ] ^ i_code[ 20 ] ^ i_code[ 21 ] ^ i_code[ 22 ] ^ i_code[ 23 ] ^ i_code[ 28 ] ^ i_code[ 29 ] ^ i_code[ 30 ] ^ i_code[ 31 ] ^ i_code[ 36 ] ^ i_code[ 37 ] ^ i_code[ 38 ];
assign o_syndrome[ 3 ] = i_code[ 8 ] ^ i_code[ 9 ] ^ i_code[ 10 ] ^ i_code[ 11 ] ^ i_code[ 12 ] ^ i_code[ 13 ] ^ i_code[ 14 ] ^ i_code[ 15 ] ^ i_code[ 24 ] ^ i_code[ 25 ] ^ i_code[ 26 ] ^ i_code[ 27 ] ^ i_code[ 28 ] ^ i_code[ 29 ] ^ i_code[ 30 ] ^ i_code[ 31 ];
assign o_syndrome[ 4 ] = i_code[ 16 ] ^ i_code[ 17 ] ^ i_code[ 18 ] ^ i_code[ 19 ] ^ i_code[ 20 ] ^ i_code[ 21 ] ^ i_code[ 22 ] ^ i_code[ 23 ] ^ i_code[ 24 ] ^ i_code[ 25 ] ^ i_code[ 26 ] ^ i_code[ 27 ] ^ i_code[ 28 ] ^ i_code[ 29 ] ^ i_code[ 30 ] ^ i_code[ 31 ];
assign o_syndrome[ 5 ] = i_code[ 32 ] ^ i_code[ 33 ] ^ i_code[ 34 ] ^ i_code[ 35 ] ^ i_code[ 36 ] ^ i_code[ 37 ] ^ i_code[ 38 ];

// Decision logic
assign o_int_sec  = parity0;
assign o_int_ded  = !parity0 && (|o_syndrome);
assign correct_bit[ 1 ] = (o_syndrome == 6'd1);
assign correct_bit[ 2 ] = (o_syndrome == 6'd2);
assign correct_bit[ 3 ] = (o_syndrome == 6'd3);
assign correct_bit[ 4 ] = (o_syndrome == 6'd4);
assign correct_bit[ 5 ] = (o_syndrome == 6'd5);
assign correct_bit[ 6 ] = (o_syndrome == 6'd6);
assign correct_bit[ 7 ] = (o_syndrome == 6'd7);
assign correct_bit[ 8 ] = (o_syndrome == 6'd8);
assign correct_bit[ 9 ] = (o_syndrome == 6'd9);
assign correct_bit[ 10 ] = (o_syndrome == 6'd10);
assign correct_bit[ 11 ] = (o_syndrome == 6'd11);
assign correct_bit[ 12 ] = (o_syndrome == 6'd12);
assign correct_bit[ 13 ] = (o_syndrome == 6'd13);
assign correct_bit[ 14 ] = (o_syndrome == 6'd14);
assign correct_bit[ 15 ] = (o_syndrome == 6'd15);
assign correct_bit[ 16 ] = (o_syndrome == 6'd16);
assign correct_bit[ 17 ] = (o_syndrome == 6'd17);
assign correct_bit[ 18 ] = (o_syndrome == 6'd18);
assign correct_bit[ 19 ] = (o_syndrome == 6'd19);
assign correct_bit[ 20 ] = (o_syndrome == 6'd20);
assign correct_bit[ 21 ] = (o_syndrome == 6'd21);
assign correct_bit[ 22 ] = (o_syndrome == 6'd22);
assign correct_bit[ 23 ] = (o_syndrome == 6'd23);
assign correct_bit[ 24 ] = (o_syndrome == 6'd24);
assign correct_bit[ 25 ] = (o_syndrome == 6'd25);
assign correct_bit[ 26 ] = (o_syndrome == 6'd26);
assign correct_bit[ 27 ] = (o_syndrome == 6'd27);
assign correct_bit[ 28 ] = (o_syndrome == 6'd28);
assign correct_bit[ 29 ] = (o_syndrome == 6'd29);
assign correct_bit[ 30 ] = (o_syndrome == 6'd30);
assign correct_bit[ 31 ] = (o_syndrome == 6'd31);
assign correct_bit[ 32 ] = (o_syndrome == 6'd32);
assign correct_bit[ 33 ] = (o_syndrome == 6'd33);
assign correct_bit[ 34 ] = (o_syndrome == 6'd34);
assign correct_bit[ 35 ] = (o_syndrome == 6'd35);
assign correct_bit[ 36 ] = (o_syndrome == 6'd36);
assign correct_bit[ 37 ] = (o_syndrome == 6'd37);
assign correct_bit[ 38 ] = (o_syndrome == 6'd38);

// Extract data bits
assign o_data[ 0 ] = correct_bit[ 3 ]? ~i_code[ 3 ] : i_code[ 3 ];
assign o_data[ 1 ] = correct_bit[ 5 ]? ~i_code[ 5 ] : i_code[ 5 ];
assign o_data[ 2 ] = correct_bit[ 6 ]? ~i_code[ 6 ] : i_code[ 6 ];
assign o_data[ 3 ] = correct_bit[ 7 ]? ~i_code[ 7 ] : i_code[ 7 ];
assign o_data[ 4 ] = correct_bit[ 9 ]? ~i_code[ 9 ] : i_code[ 9 ];
assign o_data[ 5 ] = correct_bit[ 10 ]? ~i_code[ 10 ] : i_code[ 10 ];
assign o_data[ 6 ] = correct_bit[ 11 ]? ~i_code[ 11 ] : i_code[ 11 ];
assign o_data[ 7 ] = correct_bit[ 12 ]? ~i_code[ 12 ] : i_code[ 12 ];
assign o_data[ 8 ] = correct_bit[ 13 ]? ~i_code[ 13 ] : i_code[ 13 ];
assign o_data[ 9 ] = correct_bit[ 14 ]? ~i_code[ 14 ] : i_code[ 14 ];
assign o_data[ 10 ] = correct_bit[ 15 ]? ~i_code[ 15 ] : i_code[ 15 ];
assign o_data[ 11 ] = correct_bit[ 17 ]? ~i_code[ 17 ] : i_code[ 17 ];
assign o_data[ 12 ] = correct_bit[ 18 ]? ~i_code[ 18 ] : i_code[ 18 ];
assign o_data[ 13 ] = correct_bit[ 19 ]? ~i_code[ 19 ] : i_code[ 19 ];
assign o_data[ 14 ] = correct_bit[ 20 ]? ~i_code[ 20 ] : i_code[ 20 ];
assign o_data[ 15 ] = correct_bit[ 21 ]? ~i_code[ 21 ] : i_code[ 21 ];
assign o_data[ 16 ] = correct_bit[ 22 ]? ~i_code[ 22 ] : i_code[ 22 ];
assign o_data[ 17 ] = correct_bit[ 23 ]? ~i_code[ 23 ] : i_code[ 23 ];
assign o_data[ 18 ] = correct_bit[ 24 ]? ~i_code[ 24 ] : i_code[ 24 ];
assign o_data[ 19 ] = correct_bit[ 25 ]? ~i_code[ 25 ] : i_code[ 25 ];
assign o_data[ 20 ] = correct_bit[ 26 ]? ~i_code[ 26 ] : i_code[ 26 ];
assign o_data[ 21 ] = correct_bit[ 27 ]? ~i_code[ 27 ] : i_code[ 27 ];
assign o_data[ 22 ] = correct_bit[ 28 ]? ~i_code[ 28 ] : i_code[ 28 ];
assign o_data[ 23 ] = correct_bit[ 29 ]? ~i_code[ 29 ] : i_code[ 29 ];
assign o_data[ 24 ] = correct_bit[ 30 ]? ~i_code[ 30 ] : i_code[ 30 ];
assign o_data[ 25 ] = correct_bit[ 31 ]? ~i_code[ 31 ] : i_code[ 31 ];
assign o_data[ 26 ] = correct_bit[ 33 ]? ~i_code[ 33 ] : i_code[ 33 ];
assign o_data[ 27 ] = correct_bit[ 34 ]? ~i_code[ 34 ] : i_code[ 34 ];
assign o_data[ 28 ] = correct_bit[ 35 ]? ~i_code[ 35 ] : i_code[ 35 ];
assign o_data[ 29 ] = correct_bit[ 36 ]? ~i_code[ 36 ] : i_code[ 36 ];
assign o_data[ 30 ] = correct_bit[ 37 ]? ~i_code[ 37 ] : i_code[ 37 ];
assign o_data[ 31 ] = correct_bit[ 38 ]? ~i_code[ 38 ] : i_code[ 38 ];

endmodule

